//----------------------------------------------------------------------
//  Butterfly: Add/Sub and Scaling
//----------------------------------------------------------------------
module Butterfly #(
    parameter   int WIDTH = 16,
    parameter   bit RH = 0  //  Round Half Up
)(
    input   logic signed  [WIDTH-1:0] x0_re,  //  Input Data #0 (Real)
    input   logic signed  [WIDTH-1:0] x0_im,  //  Input Data #0 (Imag)
    input   logic signed  [WIDTH-1:0] x1_re,  //  Input Data #1 (Real)
    input   logic signed  [WIDTH-1:0] x1_im,  //  Input Data #1 (Imag)
    output  logic signed  [WIDTH-1:0] y0_re,  //  Output Data #0 (Real)
    output  logic signed  [WIDTH-1:0] y0_im,  //  Output Data #0 (Imag)
    output  logic signed  [WIDTH-1:0] y1_re,  //  Output Data #1 (Real)
    output  logic signed  [WIDTH-1:0] y1_im   //  Output Data #1 (Imag)
);

logic signed [WIDTH:0]   add_re, add_im, sub_re, sub_im;

//  Add/Sub
assign  add_re = x0_re + x1_re;
assign  add_im = x0_im + x1_im;
assign  sub_re = x0_re - x1_re;
assign  sub_im = x0_im - x1_im;

//  Scaling
assign  y0_re = (add_re + RH) >>> 1;
assign  y0_im = (add_im + RH) >>> 1;
assign  y1_re = (sub_re + RH) >>> 1;
assign  y1_im = (sub_im + RH) >>> 1;

endmodule